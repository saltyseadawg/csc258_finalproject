player module(seq, check, seq_counter, playerEN, checkEN);
	input [17:0] seq;
	input [5:0] seq_counter;
	input playerEN, checkEN;
	
	output reg check;
	
	
	
endmodule;